----------------------------------------------------------------------------------
-- Engineer: Chewepe Tsate
-- 
-- Create Date: 23.10.2020 15:02:34
-- Design Name: Blowfish
-- Module Name: BlowfishHeader - Header
-- Project Name: CryptographyAlgorithms
-- Target Devices: ARM MPS2+ FPGA Prototyping Board
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package BlowfishHeader2 is

--Types
--type keyarray is array (0 to 13) of std_logic_vector(31 downto 0); --55 lots of 8 which makes 448 bits OR 13 lots of 32
type Pkeys is array (0 to 17) of std_logic_vector(31 downto 0); 
type Sboxes is array (0 to 255) of std_logic_vector(31 downto 0);
type KEYS is array (0 to 7) of std_logic_vector(31 downto 0);

--Constants
constant INITIAL_P : Pkeys := (x"243F6A88", x"85A308D3", x"13198A2E", x"03707344",
                                x"A4093822", x"299F31D0", x"082EFA98", x"EC4E6C89",
                                x"452821E6", x"38D01377", x"BE5466CF", x"34E90C6C",
                                x"C0AC29B7", x"C97C50DD", x"3F84D5B5", x"B5470917",
                                x"9216D5D9", x"8979FB1B");

constant INITAL_S0 : Sboxes := (
   x"D1310BA6",x"98DFB5AC",x"2FFD72DB",x"D01ADFB7",x"B8E1AFED",x"6A267E96",x"BA7C9045",x"F12C7F99",
   x"24A19947",x"B3916CF7",x"0801F2E2",x"858EFC16",x"636920D8",x"71574E69",x"A458FEA3",x"F4933D7E",
   x"0D95748F",x"728EB658",x"718BCD58",x"82154AEE",x"7B54A41D",x"C25A59B5",x"9C30D539",x"2AF26013",
   x"C5D1B023",x"286085F0",x"CA417918",x"B8DB38EF",x"8E79DCB0",x"603A180E",x"6C9E0E8B",x"B01E8A3E",
   x"D71577C1",x"BD314B27",x"78AF2FDA",x"55605C60",x"E65525F3",x"AA55AB94",x"57489862",x"63E81440",
   x"55CA396A",x"2AAB10B6",x"B4CC5C34",x"1141E8CE",x"A15486AF",x"7C72E993",x"B3EE1411",x"636FBC2A",
   x"2BA9C55D",x"741831F6",x"CE5C3E16",x"9B87931E",x"AFD6BA33",x"6C24CF5C",x"7A325381",x"28958677",
   x"3B8F4898",x"6B4BB9AF",x"C4BFE81B",x"66282193",x"61D809CC",x"FB21A991",x"487CAC60",x"5DEC8032",
   x"EF845D5D",x"E98575B1",x"DC262302",x"EB651B88",x"23893E81",x"D396ACC5",x"0F6D6FF3",x"83F44239",
   x"2E0B4482",x"A4842004",x"69C8F04A",x"9E1F9B5E",x"21C66842",x"F6E96C9A",x"670C9C61",x"ABD388F0",
   x"6A51A0D2",x"D8542F68",x"960FA728",x"AB5133A3",x"6EEF0B6C",x"137A3BE4",x"BA3BF050",x"7EFB2A98",
   x"A1F1651D",x"39AF0176",x"66CA593E",x"82430E88",x"8CEE8619",x"456F9FB4",x"7D84A5C3",x"3B8B5EBE",
   x"E06F75D8",x"85C12073",x"401A449F",x"56C16AA6",x"4ED3AA62",x"363F7706",x"1BFEDF72",x"429B023D",
   x"37D0D724",x"D00A1248",x"DB0FEAD3",x"49F1C09B",x"075372C9",x"80991B7B",x"25D479D8",x"F6E8DEF7",
   x"E3FE501A",x"B6794C3B",x"976CE0BD",x"04C006BA",x"C1A94FB6",x"409F60C4",x"5E5C9EC2",x"196A2463",
   x"68FB6FAF",x"3E6C53B5",x"1339B2EB",x"3B52EC6F",x"6DFC511F",x"9B30952C",x"CC814544",x"AF5EBD09",
   x"BEE3D004",x"DE334AFD",x"660F2807",x"192E4BB3",x"C0CBA857",x"45C8740F",x"D20B5F39",x"B9D3FBDB",
   x"5579C0BD",x"1A60320A",x"D6A100C6",x"402C7279",x"679F25FE",x"FB1FA3CC",x"8EA5E9F8",x"DB3222F8",
   x"3C7516DF",x"FD616B15",x"2F501EC8",x"AD0552AB",x"323DB5FA",x"FD238760",x"53317B48",x"3E00DF82",
   x"9E5C57BB",x"CA6F8CA0",x"1A87562E",x"DF1769DB",x"D542A8F6",x"287EFFC3",x"AC6732C6",x"8C4F5573",
   x"695B27B0",x"BBCA58C8",x"E1FFA35D",x"B8F011A0",x"10FA3D98",x"FD2183B8",x"4AFCB56C",x"2DD1D35B",
   x"9A53E479",x"B6F84565",x"D28E49BC",x"4BFB9790",x"E1DDF2DA",x"A4CB7E33",x"62FB1341",x"CEE4C6E8",
   x"EF20CADA",x"36774C01",x"D07E9EFE",x"2BF11FB4",x"95DBDA4D",x"AE909198",x"EAAD8E71",x"6B93D5A0",
   x"D08ED1D0",x"AFC725E0",x"8E3C5B2F",x"8E7594B7",x"8FF6E2FB",x"F2122B64",x"8888B812",x"900DF01C",
   x"4FAD5EA0",x"688FC31C",x"D1CFF191",x"B3A8C1AD",x"2F2F2218",x"BE0E1777",x"EA752DFE",x"8B021FA1",
   x"E5A0CC0F",x"B56F74E8",x"18ACF3D6",x"CE89E299",x"B4A84FE0",x"FD13E0B7",x"7CC43B81",x"D2ADA8D9",
   x"165FA266",x"80957705",x"93CC7314",x"211A1477",x"E6AD2065",x"77B5FA86",x"C75442F5",x"FB9D35CF",
   x"EBCDAF0C",x"7B3E89A0",x"D6411BD3",x"AE1E7E49",x"00250E2D",x"2071B35E",x"226800BB",x"57B8E0AF",
   x"2464369B",x"F009B91E",x"5563911D",x"59DFA6AA",x"78C14389",x"D95A537F",x"207D5BA2",x"02E5B9C5",
   x"83260376",x"6295CFA9",x"11C81968",x"4E734A41",x"B3472DCA",x"7B14A94A",x"1B510052",x"9A532915",
   x"D60F573F",x"BC9BC6E4",x"2B60A476",x"81E67400",x"08BA6FB5",x"571BE91F",x"F296EC6B",x"2A0DD915",
   x"B6636521",x"E7B9F9B6",x"FF34052E",x"C5855664",x"53B02D5D",x"A99F8FA1",x"08BA4799",x"6E85076A");

constant INITAL_S1 : Sboxes := (x"4B7A70E9",x"B5B32944",x"DB75092E",x"C4192623",x"AD6EA6B0",x"49A7DF7D",x"9CEE60B8",x"8FEDB266",
   x"ECAA8C71",x"699A17FF",x"5664526C",x"C2B19EE1",x"193602A5",x"75094C29",x"A0591340",x"E4183A3E",
   x"3F54989A",x"5B429D65",x"6B8FE4D6",x"99F73FD6",x"A1D29C07",x"EFE830F5",x"4D2D38E6",x"F0255DC1",
   x"4CDD2086",x"8470EB26",x"6382E9C6",x"021ECC5E",x"09686B3F",x"3EBAEFC9",x"3C971814",x"6B6A70A1",
   x"687F3584",x"52A0E286",x"B79C5305",x"AA500737",x"3E07841C",x"7FDEAE5C",x"8E7D44EC",x"5716F2B8",
   x"B03ADA37",x"F0500C0D",x"F01C1F04",x"0200B3FF",x"AE0CF51A",x"3CB574B2",x"25837A58",x"DC0921BD",
   x"D19113F9",x"7CA92FF6",x"94324773",x"22F54701",x"3AE5E581",x"37C2DADC",x"C8B57634",x"9AF3DDA7",
   x"A9446146",x"0FD0030E",x"ECC8C73E",x"A4751E41",x"E238CD99",x"3BEA0E2F",x"3280BBA1",x"183EB331",
   x"4E548B38",x"4F6DB908",x"6F420D03",x"F60A04BF",x"2CB81290",x"24977C79",x"5679B072",x"BCAF89AF",
   x"DE9A771F",x"D9930810",x"B38BAE12",x"DCCF3F2E",x"5512721F",x"2E6B7124",x"501ADDE6",x"9F84CD87",
   x"7A584718",x"7408DA17",x"BC9F9ABC",x"E94B7D8C",x"EC7AEC3A",x"DB851DFA",x"63094366",x"C464C3D2",
   x"EF1C1847",x"3215D908",x"DD433B37",x"24C2BA16",x"12A14D43",x"2A65C451",x"50940002",x"133AE4DD",
   x"71DFF89E",x"10314E55",x"81AC77D6",x"5F11199B",x"043556F1",x"D7A3C76B",x"3C11183B",x"5924A509",
   x"F28FE6ED",x"97F1FBFA",x"9EBABF2C",x"1E153C6E",x"86E34570",x"EAE96FB1",x"860E5E0A",x"5A3E2AB3",
   x"771FE71C",x"4E3D06FA",x"2965DCB9",x"99E71D0F",x"803E89D6",x"5266C825",x"2E4CC978",x"9C10B36A",
   x"C6150EBA",x"94E2EA78",x"A5FC3C53",x"1E0A2DF4",x"F2F74EA7",x"361D2B3D",x"1939260F",x"19C27960",
   x"5223A708",x"F71312B6",x"EBADFE6E",x"EAC31F66",x"E3BC4595",x"A67BC883",x"B17F37D1",x"018CFF28",
   x"C332DDEF",x"BE6C5AA5",x"65582185",x"68AB9802",x"EECEA50F",x"DB2F953B",x"2AEF7DAD",x"5B6E2F84",
   x"1521B628",x"29076170",x"ECDD4775",x"619F1510",x"13CCA830",x"EB61BD96",x"0334FE1E",x"AA0363CF",
   x"B5735C90",x"4C70A239",x"D59E9E0B",x"CBAADE14",x"EECC86BC",x"60622CA7",x"9CAB5CAB",x"B2F3846E",
   x"648B1EAF",x"19BDF0CA",x"A02369B9",x"655ABB50",x"40685A32",x"3C2AB4B3",x"319EE9D5",x"C021B8F7",
   x"9B540B19",x"875FA099",x"95F7997E",x"623D7DA8",x"F837889A",x"97E32D77",x"11ED935F",x"16681281",
   x"0E358829",x"C7E61FD6",x"96DEDFA1",x"7858BA99",x"57F584A5",x"1B227263",x"9B83C3FF",x"1AC24696",
   x"CDB30AEB",x"532E3054",x"8FD948E4",x"6DBC3128",x"58EBF2EF",x"34C6FFEA",x"FE28ED61",x"EE7C3C73",
   x"5D4A14D9",x"E864B7E3",x"42105D14",x"203E13E0",x"45EEE2B6",x"A3AAABEA",x"DB6C4F15",x"FACB4FD0",
   x"C742F442",x"EF6ABBB5",x"654F3B1D",x"41CD2105",x"D81E799E",x"86854DC7",x"E44B476A",x"3D816250",
   x"CF62A1F2",x"5B8D2646",x"FC8883A0",x"C1C7B6A3",x"7F1524C3",x"69CB7492",x"47848A0B",x"5692B285",
   x"095BBF00",x"AD19489D",x"1462B174",x"23820E00",x"58428D2A",x"0C55F5EA",x"1DADF43E",x"233F7061",
   x"3372F092",x"8D937E41",x"D65FECF1",x"6C223BDB",x"7CDE3759",x"CBEE7460",x"4085F2A7",x"CE77326E",
   x"A6078084",x"19F8509E",x"E8EFD855",x"61D99735",x"A969A7AA",x"C50C06C2",x"5A04ABFC",x"800BCADC",
   x"9E447A2E",x"C3453484",x"FDD56705",x"0E1E9EC9",x"DB73DBD3",x"105588CD",x"675FDA79",x"E3674340",
   x"C5C43465",x"713E38D8",x"3D28F89E",x"F16DFF20",x"153E21E7",x"8FB03D4A",x"E6E39F2B",x"DB83ADF7");

constant INITAL_S2 : Sboxes := (x"E93D5A68",x"948140F7",x"F64C261C",x"94692934",x"411520F7",x"7602D4F7",x"BCF46B2E",x"D4A20068",
   x"D4082471",x"3320F46A",x"43B7D4B7",x"500061AF",x"1E39F62E",x"97244546",x"14214F74",x"BF8B8840",
   x"4D95FC1D",x"96B591AF",x"70F4DDD3",x"66A02F45",x"BFBC09EC",x"03BD9785",x"7FAC6DD0",x"31CB8504",
   x"96EB27B3",x"55FD3941",x"DA2547E6",x"ABCA0A9A",x"28507825",x"530429F4",x"0A2C86DA",x"E9B66DFB",
   x"68DC1462",x"D7486900",x"680EC0A4",x"27A18DEE",x"4F3FFEA2",x"E887AD8C",x"B58CE006",x"7AF4D6B6",
   x"AACE1E7C",x"D3375FEC",x"CE78A399",x"406B2A42",x"20FE9E35",x"D9F385B9",x"EE39D7AB",x"3B124E8B",
   x"1DC9FAF7",x"4B6D1856",x"26A36631",x"EAE397B2",x"3A6EFA74",x"DD5B4332",x"6841E7F7",x"CA7820FB",
   x"FB0AF54E",x"D8FEB397",x"454056AC",x"BA489527",x"55533A3A",x"20838D87",x"FE6BA9B7",x"D096954B",
   x"55A867BC",x"A1159A58",x"CCA92963",x"99E1DB33",x"A62A4A56",x"3F3125F9",x"5EF47E1C",x"9029317C",
   x"FDF8E802",x"04272F70",x"80BB155C",x"05282CE3",x"95C11548",x"E4C66D22",x"48C1133F",x"C70F86DC",
   x"07F9C9EE",x"41041F0F",x"404779A4",x"5D886E17",x"325F51EB",x"D59BC0D1",x"F2BCC18F",x"41113564",
   x"257B7834",x"602A9C60",x"DFF8E8A3",x"1F636C1B",x"0E12B4C2",x"02E1329E",x"AF664FD1",x"CAD18115",
   x"6B2395E0",x"333E92E1",x"3B240B62",x"EEBEB922",x"85B2A20E",x"E6BA0D99",x"DE720C8C",x"2DA2F728",
   x"D0127845",x"95B794FD",x"647D0862",x"E7CCF5F0",x"5449A36F",x"877D48FA",x"C39DFD27",x"F33E8D1E",
   x"0A476341",x"992EFF74",x"3A6F6EAB",x"F4F8FD37",x"A812DC60",x"A1EBDDF8",x"991BE14C",x"DB6E6B0D",
   x"C67B5510",x"6D672C37",x"2765D43B",x"DCD0E804",x"F1290DC7",x"CC00FFA3",x"B5390F92",x"690FED0B",
   x"667B9FFB",x"CEDB7D9C",x"A091CF0B",x"D9155EA3",x"BB132F88",x"515BAD24",x"7B9479BF",x"763BD6EB",
   x"37392EB3",x"CC115979",x"8026E297",x"F42E312D",x"6842ADA7",x"C66A2B3B",x"12754CCC",x"782EF11C",
   x"6A124237",x"B79251E7",x"06A1BBE6",x"4BFB6350",x"1A6B1018",x"11CAEDFA",x"3D25BDD8",x"E2E1C3C9",
   x"44421659",x"0A121386",x"D90CEC6E",x"D5ABEA2A",x"64AF674E",x"DA86A85F",x"BEBFE988",x"64E4C3FE",
   x"9DBC8057",x"F0F7C086",x"60787BF8",x"6003604D",x"D1FD8346",x"F6381FB0",x"7745AE04",x"D736FCCC",
   x"83426B33",x"F01EAB71",x"B0804187",x"3C005E5F",x"77A057BE",x"BDE8AE24",x"55464299",x"BF582E61",
   x"4E58F48F",x"F2DDFDA2",x"F474EF38",x"8789BDC2",x"5366F9C3",x"C8B38E74",x"B475F255",x"46FCD9B9",
   x"7AEB2661",x"8B1DDF84",x"846A0E79",x"915F95E2",x"466E598E",x"20B45770",x"8CD55591",x"C902DE4C",
   x"B90BACE1",x"BB8205D0",x"11A86248",x"7574A99E",x"B77F19B6",x"E0A9DC09",x"662D09A1",x"C4324633",
   x"E85A1F02",x"09F0BE8C",x"4A99A025",x"1D6EFE10",x"1AB93D1D",x"0BA5A4DF",x"A186F20F",x"2868F169",
   x"DCB7DA83",x"573906FE",x"A1E2CE9B",x"4FCD7F52",x"50115E01",x"A70683FA",x"A002B5C4",x"0DE6D027",
   x"9AF88C27",x"773F8641",x"C3604C06",x"61A806B5",x"F0177A28",x"C0F586E0",x"006058AA",x"30DC7D62",
   x"11E69ED7",x"2338EA63",x"53C2DD94",x"C2C21634",x"BBCBEE56",x"90BCB6DE",x"EBFC7DA1",x"CE591D76",
   x"6F05E409",x"4B7C0188",x"39720A3D",x"7C927C24",x"86E3725F",x"724D9DB9",x"1AC15BB4",x"D39EB8FC",
   x"ED545578",x"08FCA5B5",x"D83D7CD3",x"4DAD0FC4",x"1E50EF5E",x"B161E6F8",x"A28514D9",x"6C51133C",
   x"6FD5C7E7",x"56E14EC4",x"362ABFCE",x"DDC6C837",x"D79A3234",x"92638212",x"670EFA8E",x"406000E0");

constant INITAL_S3 : Sboxes :=  (x"3A39CE37",x"D3FAF5CF",x"ABC27737",x"5AC52D1B",x"5CB0679E",x"4FA33742",x"D3822740",x"99BC9BBE",
   x"D5118E9D",x"BF0F7315",x"D62D1C7E",x"C700C47B",x"B78C1B6B",x"21A19045",x"B26EB1BE",x"6A366EB4",
   x"5748AB2F",x"BC946E79",x"C6A376D2",x"6549C2C8",x"530FF8EE",x"468DDE7D",x"D5730A1D",x"4CD04DC6",
   x"2939BBDB",x"A9BA4650",x"AC9526E8",x"BE5EE304",x"A1FAD5F0",x"6A2D519A",x"63EF8CE2",x"9A86EE22",
   x"C089C2B8",x"43242EF6",x"A51E03AA",x"9CF2D0A4",x"83C061BA",x"9BE96A4D",x"8FE51550",x"BA645BD6",
   x"2826A2F9",x"A73A3AE1",x"4BA99586",x"EF5562E9",x"C72FEFD3",x"F752F7DA",x"3F046F69",x"77FA0A59",
   x"80E4A915",x"87B08601",x"9B09E6AD",x"3B3EE593",x"E990FD5A",x"9E34D797",x"2CF0B7D9",x"022B8B51",
   x"96D5AC3A",x"017DA67D",x"D1CF3ED6",x"7C7D2D28",x"1F9F25CF",x"ADF2B89B",x"5AD6B472",x"5A88F54C",
   x"E029AC71",x"E019A5E6",x"47B0ACFD",x"ED93FA9B",x"E8D3C48D",x"283B57CC",x"F8D56629",x"79132E28",
   x"785F0191",x"ED756055",x"F7960E44",x"E3D35E8C",x"15056DD4",x"88F46DBA",x"03A16125",x"0564F0BD",
   x"C3EB9E15",x"3C9057A2",x"97271AEC",x"A93A072A",x"1B3F6D9B",x"1E6321F5",x"F59C66FB",x"26DCF319",
   x"7533D928",x"B155FDF5",x"03563482",x"8ABA3CBB",x"28517711",x"C20AD9F8",x"ABCC5167",x"CCAD925F",
   x"4DE81751",x"3830DC8E",x"379D5862",x"9320F991",x"EA7A90C2",x"FB3E7BCE",x"5121CE64",x"774FBE32",
   x"A8B6E37E",x"C3293D46",x"48DE5369",x"6413E680",x"A2AE0810",x"DD6DB224",x"69852DFD",x"09072166",
   x"B39A460A",x"6445C0DD",x"586CDECF",x"1C20C8AE",x"5BBEF7DD",x"1B588D40",x"CCD2017F",x"6BB4E3BB",
   x"DDA26A7E",x"3A59FF45",x"3E350A44",x"BCB4CDD5",x"72EACEA8",x"FA6484BB",x"8D6612AE",x"BF3C6F47",
   x"D29BE463",x"542F5D9E",x"AEC2771B",x"F64E6370",x"740E0D8D",x"E75B1357",x"F8721671",x"AF537D5D",
   x"4040CB08",x"4EB4E2CC",x"34D2466A",x"0115AF84",x"E1B00428",x"95983A1D",x"06B89FB4",x"CE6EA048",
   x"6F3F3B82",x"3520AB82",x"011A1D4B",x"277227F8",x"611560B1",x"E7933FDC",x"BB3A792B",x"344525BD",
   x"A08839E1",x"51CE794B",x"2F32C9B7",x"A01FBAC9",x"E01CC87E",x"BCC7D1F6",x"CF0111C3",x"A1E8AAC7",
   x"1A908749",x"D44FBD9A",x"D0DADECB",x"D50ADA38",x"0339C32A",x"C6913667",x"8DF9317C",x"E0B12B4F",
   x"F79E59B7",x"43F5BB3A",x"F2D519FF",x"27D9459C",x"BF97222C",x"15E6FC2A",x"0F91FC71",x"9B941525",
   x"FAE59361",x"CEB69CEB",x"C2A86459",x"12BAA8D1",x"B6C1075E",x"E3056A0C",x"10D25065",x"CB03A442",
   x"E0EC6E0E",x"1698DB3B",x"4C98A0BE",x"3278E964",x"9F1F9532",x"E0D392DF",x"D3A0342B",x"8971F21E",
   x"1B0A7441",x"4BA3348C",x"C5BE7120",x"C37632D8",x"DF359F8D",x"9B992F2E",x"E60B6F47",x"0FE3F11D",
   x"E54CDA54",x"1EDAD891",x"CE6279CF",x"CD3E7E6F",x"1618B166",x"FD2C1D05",x"848FD2C5",x"F6FB2299",
   x"F523F357",x"A6327623",x"93A83531",x"56CCCD02",x"ACF08162",x"5A75EBB5",x"6E163697",x"88D273CC",
   x"DE966292",x"81B949D0",x"4C50901B",x"71C65614",x"E6C6C7BD",x"327A140A",x"45E1D006",x"C3F27B9A",
   x"C9AA53FD",x"62A80F00",x"BB25BFE2",x"35BDD2F6",x"71126905",x"B2040222",x"B6CBCF7C",x"CD769C2B",
   x"53113EC0",x"1640E3D3",x"38ABBD60",x"2547ADF0",x"BA38209C",x"F746CE76",x"77AFA1C5",x"20756060",
   x"85CBFE4E",x"8AE88DD8",x"7AAAF9B0",x"4CF9AA7E",x"1948C25C",x"02FB8A8C",x"01C36AE4",x"D6EBE1F9",
   x"90D4F869",x"A65CDEA0",x"3F09252D",x"C208E69F",x"B74E6132",x"CE77E25B",x"578FDFE3",x"3AC372E6");

end;